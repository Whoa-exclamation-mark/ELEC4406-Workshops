library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
  
  
entity blank_entity is
end blank_entity;
	
	
architecture blank_entity_rtl of blank_entity is 

begin 
	
end blank_entity_rtl;